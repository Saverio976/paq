module paq
